`timescale 1ns/1ns
module ArrayConvLayerCtrl_tb#(parameter
    num_pe_row = 16,
    num_pe_col = 16,
    total_num_pe = num_pe_row * num_pe_col,
    //parameter for conv layer controller
    max_outch_per_time = 256,
    ACCFIFO_size = 32,
    tiled_col_size = ACCFIFO_size,
    inch_group_size = 16,
    outch_group_size = (max_outch_per_time + num_pe_col - 1) / num_pe_col,
    //parameters for PE and FoFIR
	nb_taps = 11,
	activation_width = 16,
	compressed_act_width = activation_width + 1,
	weight_width = 16,
	tap_width = 24,
	weight_bpr_width = ((weight_width+1)/2)*3,
	act_bpr_width = ((activation_width+1)/2)*3,
	ETC_width = 4,
	width_current_tap = nb_taps > 8 ? 4 : 3,
	output_width = tap_width
    )();
    /**** Ports from conv_one_row_ctrl to control the PE array (started with ``pe_ctrl/data")*****/
    // AFIFO data
        logic [num_pe_row-1: 0][compressed_act_width-1: 0] pe_data_compressed_act_in;
        logic [num_pe_col-1: 0][compressed_act_width-1: 0] pe_data_last_row_shadow_AFIFO_data_in;
    // configuration
        logic [total_num_pe-1: 0][4-1: 0] pe_ctrl_n_ap;
    // control ports for PAMAC
        logic [total_num_pe-1: 0][3-1: 0] pe_ctrl_PAMAC_BPEB_sel;
        logic [total_num_pe-1: 0] pe_ctrl_PAMAC_DFF_en;
        logic [total_num_pe-1: 0] pe_ctrl_PAMAC_first_cycle;
        logic [total_num_pe-1: 0] pe_ctrl_PAMAC_MDecomp;
        logic [total_num_pe-1: 0] pe_ctrl_PAMAC_AWDecomp;
    // control ports for FoFIR
        logic [total_num_pe-1: 0][width_current_tap-1: 0] pe_ctrl_current_tap;
        logic [total_num_pe-1: 0][nb_taps-1: 0] pe_ctrl_DRegs_en;
        logic [total_num_pe-1: 0][nb_taps-1: 0] pe_ctrl_DRegs_clr;
        logic [total_num_pe-1: 0][nb_taps-1: 0] pe_ctrl_DRegs_in_sel;
        logic [total_num_pe-1: 0] pe_ctrl_index_update_en;
        logic [total_num_pe-1: 0] pe_ctrl_out_mux_sel;
        logic [total_num_pe-1: 0] pe_ctrl_out_reg_en;
    // control ports for FIFOs
        logic [total_num_pe-1: 0] pe_ctrl_AFIFO_write;
        logic [total_num_pe-1: 0] pe_ctrl_AFIFO_read; 
        logic [total_num_pe-1: 0] pe_ctrl_ACCFIFO_write;
        logic [total_num_pe-1: 0] pe_ctrl_ACCFIFO_read; //read when computing 
        logic [total_num_pe-1: 0] pe_ctrl_ACCFIFO_read_to_outbuffer;//read when let data goto out buffer
        logic [total_num_pe-1: 0] pe_ctrl_out_mux_sel_PE;// 0 is from ACCFIFO; 1 is from left PE
        logic [total_num_pe-1: 0] pe_ctrl_out_to_right_pe_en;	
        logic [total_num_pe-1: 0] pe_ctrl_add_zero;
        logic [total_num_pe-1: 0] pe_ctrl_feed_zero_to_accfifo;
        logic [total_num_pe-1: 0] pe_ctrl_accfifo_head_to_tail;
        logic [num_pe_col-1: 0] pe_ctrl_last_row_shadow_AFIFO_write;
    /**** End of Ports to control the PE array***/
    /**** Ports from PE array for some info ****/
        logic [total_num_pe-1: 0][width_current_tap-1: 0] pe_ctrl_PD0;
        logic [total_num_pe-1: 0] pe_ctrl_AFIFO_full;
        logic [total_num_pe-1: 0] pe_ctrl_AFIFO_empty;
        logic [total_num_pe-1: 0][compressed_act_width-1: 0] pe_data_afifo_out;
        logic [total_num_pe-1: 0] pe_ctrl_ACCFIFO_empty;
    /**** End of Ports from PE array for some info****/
    /**** Ports of some weights info; generated by this module*****************/
        logic [num_pe_col-1: 0][weight_width*nb_taps-1: 0] WRegs;
        logic [num_pe_col-1: 0][weight_bpr_width*nb_taps-1: 0] WBPRs;
        logic [num_pe_col-1: 0][ETC_width*nb_taps-1: 0] WETCs;
    /**** End of ports for weights info**************/
    /***** Ports from this module to schedule the whole convolutional layer***/
        logic [total_num_pe-1: 0] pe_ctrl_which_accfifo_for_compute;
        logic [total_num_pe-1: 0] pe_ctrl_compute_AFIFO_read_delay_enable;
        logic [total_num_pe-1: 0] pe_ctrl_which_afifo_for_compute;
    /******* End of Conv Layer Ctrl Ports********/
        logic array_next_cycle_data_to_outbuff_valid;
        logic clk;
        logic rst_n;
        logic [num_pe_row-1: 0][output_width-1:0] out_fr_rightest_PE_even_col;    // %2 = 0
        logic [num_pe_row-1: 0][output_width-1:0] out_fr_rightest_PE_odd_col;  
    initial begin
        clk = 0;
        forever begin
            #10 clk = ~clk;
        end
    end
    ArrayConvLayerCtrl #(
        .num_pe_col(num_pe_col),
        .num_pe_row(num_pe_row),
        .max_outch_per_time(max_outch_per_time),
        .ACCFIFO_size(ACCFIFO_size),
        .inch_group_size(inch_group_size),
        .nb_taps(nb_taps),
        .activation_width(activation_width),
        .weight_width(weight_width),
        .tap_width(tap_width),
        .ETC_width(ETC_width)
    ) DUT_Ctrl(
    	.pe_data_compressed_act_in               (pe_data_compressed_act_in               ),
        .pe_data_last_row_shadow_AFIFO_data_in   (pe_data_last_row_shadow_AFIFO_data_in   ),
        .pe_ctrl_n_ap                            (pe_ctrl_n_ap                            ),
        .pe_ctrl_PAMAC_BPEB_sel                  (pe_ctrl_PAMAC_BPEB_sel                  ),
        .pe_ctrl_PAMAC_DFF_en                    (pe_ctrl_PAMAC_DFF_en                    ),
        .pe_ctrl_PAMAC_first_cycle               (pe_ctrl_PAMAC_first_cycle               ),
        .pe_ctrl_PAMAC_MDecomp                   (pe_ctrl_PAMAC_MDecomp                   ),
        .pe_ctrl_PAMAC_AWDecomp                  (pe_ctrl_PAMAC_AWDecomp                  ),
        .pe_ctrl_current_tap                     (pe_ctrl_current_tap                     ),
        .pe_ctrl_DRegs_en                        (pe_ctrl_DRegs_en                        ),
        .pe_ctrl_DRegs_clr                       (pe_ctrl_DRegs_clr                       ),
        .pe_ctrl_DRegs_in_sel                    (pe_ctrl_DRegs_in_sel                    ),
        .pe_ctrl_index_update_en                 (pe_ctrl_index_update_en                 ),
        .pe_ctrl_out_mux_sel                     (pe_ctrl_out_mux_sel                     ),
        .pe_ctrl_out_reg_en                      (pe_ctrl_out_reg_en                      ),
        .pe_ctrl_AFIFO_write                     (pe_ctrl_AFIFO_write                     ),
        .pe_ctrl_AFIFO_read                      (pe_ctrl_AFIFO_read                      ),
        .pe_ctrl_ACCFIFO_write                   (pe_ctrl_ACCFIFO_write                   ),
        .pe_ctrl_ACCFIFO_read                    (pe_ctrl_ACCFIFO_read                    ),
        .pe_ctrl_ACCFIFO_read_to_outbuffer       (pe_ctrl_ACCFIFO_read_to_outbuffer       ),
        .pe_ctrl_out_mux_sel_PE                  (pe_ctrl_out_mux_sel_PE                  ),
        .pe_ctrl_out_to_right_pe_en              (pe_ctrl_out_to_right_pe_en              ),
        .pe_ctrl_add_zero                        (pe_ctrl_add_zero                        ),
        .pe_ctrl_feed_zero_to_accfifo            (pe_ctrl_feed_zero_to_accfifo            ),
        .pe_ctrl_accfifo_head_to_tail            (pe_ctrl_accfifo_head_to_tail            ),
        .pe_ctrl_last_row_shadow_AFIFO_write     (pe_ctrl_last_row_shadow_AFIFO_write     ),
        .pe_ctrl_PD0                             (pe_ctrl_PD0                             ),
        .pe_ctrl_AFIFO_full                      (pe_ctrl_AFIFO_full                      ),
        .pe_ctrl_AFIFO_empty                     (pe_ctrl_AFIFO_empty                     ),
        .pe_data_afifo_out                       (pe_data_afifo_out                       ),
        .pe_ctrl_ACCFIFO_empty                   (pe_ctrl_ACCFIFO_empty                   ),
        .WRegs                                   (WRegs                                   ),
        .WBPRs                                   (WBPRs                                   ),
        .WETCs                                   (WETCs                                   ),
        .pe_ctrl_which_accfifo_for_compute       (pe_ctrl_which_accfifo_for_compute       ),
        .pe_ctrl_compute_AFIFO_read_delay_enable (pe_ctrl_compute_AFIFO_read_delay_enable ),
        .pe_ctrl_which_afifo_for_compute         (pe_ctrl_which_afifo_for_compute         ),
        .array_next_cycle_data_to_outbuff_valid  (array_next_cycle_data_to_outbuff_valid  ),
        .clk                                     (clk                                     )
    );
    PEArray_for_power_analysis #(
        .num_pe_row(num_pe_row),
        .num_pe_col(num_pe_col),
        .nb_taps(nb_taps),
        .activation_width(activation_width),
        .weight_width(weight_width),
        .tap_width(tap_width),
        .ETC_width(ETC_width)
    )u_PEArray_for_power_analysis(
    	.pe_data_compressed_act_in               (pe_data_compressed_act_in               ),
        .pe_data_last_row_shadow_AFIFO_data_in   (pe_data_last_row_shadow_AFIFO_data_in   ),
        .pe_ctrl_n_ap                            (pe_ctrl_n_ap                            ),
        .pe_ctrl_PAMAC_BPEB_sel                  (pe_ctrl_PAMAC_BPEB_sel                  ),
        .pe_ctrl_PAMAC_DFF_en                    (pe_ctrl_PAMAC_DFF_en                    ),
        .pe_ctrl_PAMAC_first_cycle               (pe_ctrl_PAMAC_first_cycle               ),
        .pe_ctrl_PAMAC_MDecomp                   (pe_ctrl_PAMAC_MDecomp                   ),
        .pe_ctrl_PAMAC_AWDecomp                  (pe_ctrl_PAMAC_AWDecomp                  ),
        .pe_ctrl_current_tap                     (pe_ctrl_current_tap                     ),
        .pe_ctrl_DRegs_en                        (pe_ctrl_DRegs_en                        ),
        .pe_ctrl_DRegs_clr                       (pe_ctrl_DRegs_clr                       ),
        .pe_ctrl_DRegs_in_sel                    (pe_ctrl_DRegs_in_sel                    ),
        .pe_ctrl_index_update_en                 (pe_ctrl_index_update_en                 ),
        .pe_ctrl_out_mux_sel                     (pe_ctrl_out_mux_sel                     ),
        .pe_ctrl_out_reg_en                      (pe_ctrl_out_reg_en                      ),
        .pe_ctrl_AFIFO_write                     (pe_ctrl_AFIFO_write                     ),
        .pe_ctrl_AFIFO_read                      (pe_ctrl_AFIFO_read                      ),
        .pe_ctrl_ACCFIFO_write                   (pe_ctrl_ACCFIFO_write                   ),
        .pe_ctrl_ACCFIFO_read                    (pe_ctrl_ACCFIFO_read                    ),
        .pe_ctrl_ACCFIFO_read_to_outbuffer       (pe_ctrl_ACCFIFO_read_to_outbuffer       ),
        .pe_ctrl_out_mux_sel_PE                  (pe_ctrl_out_mux_sel_PE                  ),
        .pe_ctrl_out_to_right_pe_en              (pe_ctrl_out_to_right_pe_en              ),
        .pe_ctrl_add_zero                        (pe_ctrl_add_zero                        ),
        .pe_ctrl_feed_zero_to_accfifo            (pe_ctrl_feed_zero_to_accfifo            ),
        .pe_ctrl_accfifo_head_to_tail            (pe_ctrl_accfifo_head_to_tail            ),
        .pe_ctrl_which_accfifo_for_compute       (pe_ctrl_which_accfifo_for_compute       ),
        .pe_ctrl_which_afifo_for_compute         (pe_ctrl_which_afifo_for_compute         ),
        .pe_ctrl_compute_AFIFO_read_delay_enable (pe_ctrl_compute_AFIFO_read_delay_enable ),
        .pe_ctrl_last_row_shadow_AFIFO_write     (pe_ctrl_last_row_shadow_AFIFO_write     ),
        .pe_ctrl_PD0                             (pe_ctrl_PD0                             ),
        .pe_ctrl_AFIFO_full                      (pe_ctrl_AFIFO_full                      ),
        .pe_ctrl_AFIFO_empty                     (pe_ctrl_AFIFO_empty                     ),
        .pe_data_afifo_out                       (pe_data_afifo_out                       ),
        .WRegs                                   (WRegs                                   ),
        .WBPRs                                   (WBPRs                                   ),
        .WETCs                                   (WETCs                                   ),
        .out_fr_rightest_PE_even_col             (out_fr_rightest_PE_even_col             ),
        .out_fr_rightest_PE_odd_col              (out_fr_rightest_PE_odd_col              ),
        .pe_ctrl_ACCFIFO_empty                   (pe_ctrl_ACCFIFO_empty                   ),
        .clk                                     (clk                                     ),
        .rst_n                                   (rst_n                                   )
    );
    /************ Helper Variables********************/
    int kernel_size_per_layer[52] = '{3,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1,3,1,1};
    int is_depthwise[52] = '{0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0,1,0,0};
    int fm_size_per_layer[52] = '{226,114,112,112,114,56,56,58,56,56,58,28,28,30,28,28,30,28,28,30,14,14,16,14,14,16,14,14,16,14,14,16,14,14,16,14,14,16,14,14,16,7,7,9,7,7,9,7,7,9,7,7};
    int in_ch_per_layer[52] = '{3,32,32,16,96,96,24,144,144,24,144,144,32,192,192,32,192,192,32,192,192,64,384,384,64,384,384,64,384,384,64,384,384,96,576,576,96,576,576,96,576,576,160,960,960,160,960,960,160,960,960,320};
    int out_ch_per_layer[52] = '{32,32,16,96,96,24,144,144,24,144,144,32,192,192,32,192,192,32,192,192,64,384,384,64,384,384,64,384,384,64,384,384,96,576,576,96,576,576,96,576,576,160,960,960,160,960,960,160,960,960,320,1280};
    int stride_per_layer[52] = '{2,1,1,1,2,1,1,1,1,1,2,1,1,1,1,1,1,1,1,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,1,1,1,1,1,1,1,1,1,1,1};

    int start_layer;
    int end_layer;
    int current_layer;
    /******Main**********/
    initial begin
        string act_file_path;
        string act_dir_path;
        string weight_file_path;
        string weight_file_name;
        string weight_full_path;
        int kernel_size;
        string layer_str;
        int log_fp;
        int total_op_this_layer;
        logic [64-1: 0] start_time;
        logic [64-1: 0] end_time;
        int cycle_this_layer;
        start_layer = 1;
        end_layer = 52;
        act_dir_path = "C:/Users/jy/Desktop/mopu-testbench/testdata/mobilenet";
        weight_file_path = {act_dir_path, "/weights"};
        rst_n = 1;
        #5;
        rst_n = 0;
        #20;
        rst_n = 1;
        @(posedge clk);
        log_fp = $fopen("PerLayerCyclePerf.log", "w");
        $fdisplay(log_fp, "Layer_Index\tIsDepthwise\tInCh\tOutCh\tInfmSize\tTime\tNumberOfCycle\tPerformance(Op/Cycle)");
        for(current_layer = start_layer; current_layer<end_layer;current_layer++) begin
            start_time = $time;
            kernel_size = kernel_size_per_layer[current_layer];
            if(stride_per_layer[current_layer] != 1) begin
                continue;
            end
            $display("@%t, Start the %d-th layer.", $time, current_layer);
            layer_str.itoa(current_layer);
            act_file_path = {act_dir_path, "/act_conv_", layer_str};
            if(is_depthwise[current_layer] == 1) begin
                act_file_path = {act_file_path, "_dw"};
            end
            weight_file_name = {"conv", layer_str, "weight.dat"};
            weight_full_path = {weight_file_path, "/", weight_file_name};
            //DUT_Ctrl.load_weights_this_layer_from_file(weight_full_path, kernel_size_per_layer[current_layer]);
            if(is_depthwise[current_layer] == 1) begin
                $display("The %d-th layer is dwconv.", current_layer);
                DUT_Ctrl.dw_conv_one_layer(
                    act_file_path,
                    weight_full_path,
                    stride_per_layer[current_layer],
                    out_ch_per_layer[current_layer],
                    fm_size_per_layer[current_layer],
                    kernel_size_per_layer[current_layer]
                );
            end
            else begin
                $display("The %d-th layer is normal_conv.", current_layer);
                DUT_Ctrl.normal_conv_one_layer(
                    act_file_path,
                    weight_full_path,
                    in_ch_per_layer[current_layer],
                    out_ch_per_layer[current_layer],
                    stride_per_layer[current_layer],
                    fm_size_per_layer[current_layer],
                    kernel_size_per_layer[current_layer]
                );
                

            end
            end_time = $time;
            if(is_depthwise[current_layer] == 1) begin
                total_op_this_layer = (fm_size_per_layer[current_layer] - 2) * (fm_size_per_layer[current_layer] - 2) * out_ch_per_layer[current_layer] * kernel_size_per_layer[current_layer] * kernel_size_per_layer[current_layer];
            end
            else begin
                total_op_this_layer = fm_size_per_layer[current_layer]*fm_size_per_layer[current_layer]*out_ch_per_layer[current_layer]*kernel_size_per_layer[current_layer]*kernel_size_per_layer[current_layer]*in_ch_per_layer[current_layer];
            end
            cycle_this_layer = (end_time - start_time)/20;
            if(stride_per_layer[current_layer]==1) begin
                $fdisplay(
                    log_fp, 
                    "%d\t\t%s\t%d\t%d\t%d\t%t\t%d\t%d", 
                    current_layer, is_depthwise[current_layer]?"Yes":"No",
                    in_ch_per_layer[current_layer], out_ch_per_layer[current_layer],
                    fm_size_per_layer[current_layer], end_time-start_time,
                    cycle_this_layer, total_op_this_layer/cycle_this_layer
                );
                $display(
                    "layer_idx:%d\tDepthWise:%s\tInCh:%d\tOutCh:%d\tfmsize:%d\tElapsedTime(ns):%t\t#Cycle:%d\tOP/Cycle:%d", 
                    current_layer, is_depthwise[current_layer]?"Yes":"No",
                    in_ch_per_layer[current_layer], out_ch_per_layer[current_layer],
                    fm_size_per_layer[current_layer], end_time-start_time,
                    cycle_this_layer, total_op_this_layer/cycle_this_layer
                );
            end
            else begin
                $fdisplay(log_fp, "%d\tN/A\tN/A\tN/A\tN/A\tN/A\tN/A\tN/A", current_layer);
            end
        end
        $fclose(log_fp);
        $finish;
    end
endmodule